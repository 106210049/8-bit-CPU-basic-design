// Temporary file for syntax check
module vector;
endmodule
